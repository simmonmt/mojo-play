library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity decode is
    Port ( D_IN : in  STD_LOGIC_VECTOR (3 downto 0);
           SZ_OUT : out  STD_LOGIC_VECTOR (2 downto 0));
end decode;

architecture Behavioral of decode is

begin


end Behavioral;

